module Reg_E (clk,rst,stall,jb,pc_in,rs1_data_in,rs2_data_in,imm_in,pc_out,rs1_data_out,rs2_data_out,imm_out);
    input clk,rst,stall,jb;
    input [31:0] rs1_data_in,rs2_data_in,imm_in;
	input [15:0] pc_in;
	output reg[15:0] pc_out;
    output reg[31:0] rs1_data_out,rs2_data_out,imm_out;
    
    always @(posedge clk or posedge rst) 
    begin
        if (rst) 
        begin
            pc_out <= 16'b0;    
            rs1_data_out <=32'b0;
            rs2_data_out <= 32'b0;    
            imm_out <= 32'b0;    
        end
        else
        begin
            if (stall | jb )  //OR    ????
            begin
                pc_out <= pc_in;    
                rs1_data_out <= 32'b0;               /////    flush????
                rs2_data_out <= 32'b0;    
                imm_out <= 32'b0;   
            end
            else
            begin                
                pc_out <= pc_in;    
                rs1_data_out <= rs1_data_in;
                rs2_data_out <= rs2_data_in;    
                imm_out <= imm_in;             
            end
        end    
    end
endmodule